module robo_core (
	input clk,    // Clock
	input rst_n,  // Asynchronous reset active low
	input front,
	input left,

	output reg foward,
	output reg turn_left
);




endmodule
